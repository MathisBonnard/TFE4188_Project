cicsimgen tran

*Nothing here

.lib  "/opt/pdk/share/pdk/sky130B/libs.tech/ngspice/sky130.lib.spice" tt_mm

.lib "../../../tech/ngspice/temperature.spi" Tt

.lib "../../../tech/ngspice/supply.spi" Vt


*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
.include ../../../work/xsch/RPLY_TEMPSENS.spice

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------

*If seed needed, add "seed=4 in the option list
.option TNOM=27 GMIN=1e-15 reltol=1e-6 abstol=1e-6 keepopinfo noopiter gminsteps=5
.temp 75

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
*VDD  VDD_1V8  VSS  pwl 0 0 10n {AVDD}
VDD   VDD_1V8  VSS  dc  1.8

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
XDUT VDD_1V8 VSS Vtop Vbot Vgate RPLY_TEMPSENS

*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------

.save v(VDD_1V8) v(VSS) v(Vtop) v(Vbot) v(Vgate) v(XDUT.inpos) i(V1)

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 100p 2n 0


tran 5000p 10u
*dc temp 0 100 1

write
quit

.endc

.end

